interface intf(input bit clk, input bit rst);

	logic [width-1:0]data_in;
	logic data_ready;
	logic d_out1;

endinterface
