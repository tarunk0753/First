package my_package;
	`include"macros.svh"
	import uvm_pkg::*
	`include "my_env.svh"
	`include "my_agent.svh"
	`include "my_test.svh"

endpackage; my_pkg



