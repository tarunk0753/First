class my_component extends uvm_component;
'uvm_component_utila(my_component)

function new (string name, parent);
super.new(name, parent);
endfunction:new




