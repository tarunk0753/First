class my_transaction
`uvm_object_utils(my_transaction)

rand bit cmd; ///variables



function new (string name ="");
super.new(name);
endfunction:new

endclass: my_transaction
